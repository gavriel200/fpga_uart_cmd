module gw_gao(
    \_printer/state[1] ,
    \_printer/state[0] ,
    \state[1] ,
    \state[0] ,
    \_tx/state[1] ,
    \_tx/state[0] ,
    \_start/state[1] ,
    \_start/state[0] ,
    \_printer/enable ,
    \_tx/enable ,
    \_start/start_state[1] ,
    \_start/start_state[0] ,
    \start_state[1] ,
    \start_state[0] ,
    clk,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \_printer/state[1] ;
input \_printer/state[0] ;
input \state[1] ;
input \state[0] ;
input \_tx/state[1] ;
input \_tx/state[0] ;
input \_start/state[1] ;
input \_start/state[0] ;
input \_printer/enable ;
input \_tx/enable ;
input \_start/start_state[1] ;
input \_start/start_state[0] ;
input \start_state[1] ;
input \start_state[0] ;
input clk;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \_printer/state[1] ;
wire \_printer/state[0] ;
wire \state[1] ;
wire \state[0] ;
wire \_tx/state[1] ;
wire \_tx/state[0] ;
wire \_start/state[1] ;
wire \_start/state[0] ;
wire \_printer/enable ;
wire \_tx/enable ;
wire \_start/start_state[1] ;
wire \_start/start_state[0] ;
wire \start_state[1] ;
wire \start_state[0] ;
wire clk;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i({\_start/state[1] ,\_start/state[0] }),
    .data_i({\_printer/state[1] ,\_printer/state[0] ,\state[1] ,\state[0] ,\_tx/state[1] ,\_tx/state[0] ,\_start/state[1] ,\_start/state[0] ,\_printer/enable ,\_tx/enable ,\_start/start_state[1] ,\_start/start_state[0] ,\start_state[1] ,\start_state[0] }),
    .clk_i(clk)
);

endmodule
