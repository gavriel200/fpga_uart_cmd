module loopback(
    port_list
);

// when active just takes in rx and puts it in tx.
// need to make sure that its done before continueing with the states

    
endmodule